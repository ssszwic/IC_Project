module Tb;

endmodule
